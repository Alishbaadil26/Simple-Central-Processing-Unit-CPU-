library verilog;
use verilog.vl_types.all;
entity lab5Combined_vlg_vec_tst is
end lab5Combined_vlg_vec_tst;
